module triumph_wb_stage();





endmodule