module triumph_wb_stage(
    input  wire        clk_i,
    input  wire        rst_i
);





endmodule