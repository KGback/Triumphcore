`timescale 1ns / 1ps

module tb;

logic clk_i;
logic rstn_i;

localparam CLK_PERIOD = 20;

initial begin
    do  begin
        #(CLK_PERIOD/2) clk_i = 1;    
        #(CLK_PERIOD/2) clk_i = 0;    
    end 
    while (1);
end

initial begin
    rstn_i = 1;
    #40 rstn_i = 0;
    #40 rstn_i = 1;
    $display("===============================");
    $display("       simulation begin        ");
    $display("===============================");
    #50000;
    $finish;
end

//initial begin
//    while (1) begin
//        #20;
//      // $display("PC: 0x%x",dut.pc); 
//    end
//end
//          


triumphcore_wrapper dut(
    .clk_i              ( clk_i             ),
    .rstn_i              ( rstn_i             )
    );


endmodule
